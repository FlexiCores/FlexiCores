module tb;

endmodule : tb
