
// 	Sun Nov  8 13:13:20 2020
//	antony
//	fenrir

module core_synth (CLK, RSTN, IPORT, OPORT, PC, INSTR);

output [3:0] OPORT;
output [6:0] PC;
input CLK;
input [7:0] INSTR;
input [3:0] IPORT;
input RSTN;
wire drc_ipo_n108;
wire drc_ipo_n106;
wire drc_ipo_n104;
wire drc_ipo_n102;
wire drc_ipo_n119;
wire slo_n214;
wire drc_ipo_n100;
wire drc_ipo_n117;
wire \dpath_rf_rf7[3] ;
wire \dpath_rf_rf7[2] ;
wire \dpath_rf_rf7[1] ;
wire \dpath_rf_rf7[0] ;
wire \dpath_rf_rf6[3] ;
wire \dpath_rf_rf6[2] ;
wire \dpath_rf_rf6[1] ;
wire \dpath_rf_rf6[0] ;
wire \dpath_rf_rf5[3] ;
wire \dpath_rf_rf5[2] ;
wire \dpath_rf_rf5[1] ;
wire \dpath_rf_rf5[0] ;
wire \dpath_rf_rf4[3] ;
wire \dpath_rf_rf4[2] ;
wire \dpath_rf_rf4[1] ;
wire \dpath_rf_rf4[0] ;
wire \dpath_rf_rf3[3] ;
wire \dpath_rf_rf3[2] ;
wire \dpath_rf_rf3[1] ;
wire \dpath_rf_rf3[0] ;
wire \dpath_rf_rf2[3] ;
wire \dpath_rf_rf2[2] ;
wire \dpath_rf_rf2[1] ;
wire \dpath_rf_rf2[0] ;
wire \dpath_A[3] ;
wire \dpath_A[2] ;
wire \dpath_A[1] ;
wire \dpath_A[0] ;
wire dpath__PC_n_15;
wire dpath_n_3;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire dpath_n_2;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire dpath_n_1;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire dpath_n_0;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire dpath_rf_n_34;
wire dpath_rf_n_33;
wire dpath_rf_n_32;
wire dpath_rf_n_31;
wire n_0_83;
wire n_0_84;
wire dpath_rf_n_30;
wire dpath_rf_n_29;
wire dpath_rf_n_28;
wire dpath_rf_n_27;
wire n_0_85;
wire dpath_rf_n_26;
wire dpath_rf_n_25;
wire dpath_rf_n_24;
wire dpath_rf_n_23;
wire n_0_86;
wire n_0_87;
wire dpath_rf_n_22;
wire dpath_rf_n_21;
wire dpath_rf_n_20;
wire dpath_rf_n_19;
wire n_0_88;
wire n_0_89;
wire dpath_rf_n_18;
wire dpath_rf_n_17;
wire dpath_rf_n_16;
wire dpath_rf_n_15;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire dpath_rf_n_14;
wire dpath_rf_n_13;
wire dpath_rf_n_12;
wire dpath_rf_n_11;
wire n_0_93;
wire n_0_94;
wire dpath_rf_n_3;
wire dpath_rf_n_2;
wire dpath_rf_n_1;
wire dpath_rf_n_0;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire dpath__PC_n_7;
wire dpath__PC_n_8;
wire n_0_102;
wire dpath__PC_n_9;
wire n_0_103;
wire dpath__PC_n_10;
wire n_0_104;
wire dpath__PC_n_11;
wire n_0_105;
wire dpath__PC_n_12;
wire n_0_106;
wire dpath__PC_n_13;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire drc_ipo_n87;
wire drc_ipo_n96;
wire drc_ipo_n94;
wire drc_ipo_n90;
wire drc_ipo_n95;
wire drc_ipo_n91;
wire drc_ipo_n88;
wire drc_ipo_n98;
wire drc_ipo_n93;
wire drc_ipo_n97;
wire drc_ipo_n92;
wire drc_ipo_n86;
wire drc_ipo_n85;
wire drc_ipo_n89;
wire drc_ipo_n84;
wire drc_ipo_n83;
wire drc_ipo_n82;
wire drc_ipo_n81;
wire drc_ipo_n80;
wire drc_ipo_n79;
wire drc_ipo_n78;
wire drc_ipo_n77;
wire drc_ipo_n76;
wire drc_ipo_n75;
wire drc_ipo_n74;
wire drc_ipo_n73;
wire drc_ipo_n72;
wire drc_ipo_n71;
wire drc_ipo_n109;
wire drc_ipo_n110;
wire drc_ipo_n111;
wire drc_ipo_n112;
wire drc_ipo_n113;
wire drc_ipo_n114;
wire drc_ipo_n115;
wire drc_ipo_n120;
wire sgo___n121;
wire sgo___n122;
wire sgo__n123;
wire sgo___n124;
wire sgo___n125;
wire sgo___n126;
wire sgo___n127;
wire sgo___n_3_121;
wire sgo___n_3_122;
wire sgo___n_3_125;
wire sgo___n_3_126;
wire sgo___n_2_121;
wire sgo___n_2_122;
wire sgo___n_2_123;
wire sgo___n_2_124;
wire sgo__n_1_121;
wire sgo___n_1_123;
wire sgo___n_1_124;
wire sgo___n_1_125;
wire sgo___n_1_126;
wire sgo__n131;
wire sgo__n133;
wire slo___n135;
wire slo___n136;
wire slo___n141;
wire slo___n142;
wire slo___n149;
wire slo___n150;
wire slo___n163;
wire slo___n164;
wire slo___n190;
wire slo___n191;
wire slo___n196;
wire slo___n197;
wire slo___n204;
wire slo___n215;
wire slo___n216;
wire slo___n223;
wire slo___n224;
wire slo___n231;
wire slo___n232;


INV4 i_0_162 (.X (n_0_123), .A (PC[4]));
INV4 i_0_161 (.X (n_0_122), .A (PC[2]));
INV4 i_0_160 (.X (n_0_121), .A (PC[0]));
INV4 i_0_159 (.X (n_0_120), .A (INSTR[7]));
INV4 i_0_158 (.X (n_0_119), .A (INSTR[6]));
INV4 i_0_157 (.X (n_0_118), .A (INSTR[5]));
INV4 i_0_156 (.X (n_0_117), .A (INSTR[4]));
INV4 i_0_155 (.X (n_0_116), .A (INSTR[2]));
INV4 i_0_154 (.X (n_0_115), .A (INSTR[1]));
INV4 i_0_153 (.X (n_0_114), .A (INSTR[0]));
NAND2 i_0_152 (.X (n_0_113), .A1 (INSTR[7]), .A2 (drc_ipo_n114));
NAND2 i_0_151 (.X (n_0_112), .A1 (PC[1]), .A2 (PC[0]));
NOR2 i_0_150 (.X (n_0_111), .A1 (n_0_122), .A2 (n_0_112));
NAND2 i_0_149 (.X (n_0_110), .A1 (PC[3]), .A2 (sgo___n_3_122));
NOR2 i_0_148 (.X (n_0_109), .A1 (n_0_123), .A2 (n_0_110));
NAND2 i_0_147 (.X (n_0_108), .A1 (PC[5]), .A2 (n_0_109));
XNOR i_0_146 (.X (n_0_107), .A1 (PC[6]), .A2 (n_0_108));
MX2 i_0_145 (.X (dpath__PC_n_13), .A (INSTR[6]), .B (slo___n216), .S (drc_ipo_n82));
XOR i_0_144 (.X (n_0_106), .A1 (PC[5]), .A2 (n_0_109));
MX2 i_0_143 (.X (dpath__PC_n_12), .A (INSTR[5]), .B (slo___n142), .S (drc_ipo_n82));
XNOR i_0_142 (.X (n_0_105), .A1 (PC[4]), .A2 (n_0_110));
MX2 i_0_141 (.X (dpath__PC_n_11), .A (INSTR[4]), .B (n_0_105), .S (drc_ipo_n82));
XOR i_0_140 (.X (n_0_104), .A1 (PC[3]), .A2 (sgo___n_3_122));
MX2 i_0_139 (.X (dpath__PC_n_10), .A (INSTR[3]), .B (slo___n136), .S (drc_ipo_n82));
XNOR i_0_138 (.X (n_0_103), .A1 (PC[2]), .A2 (n_0_112));
MX2 i_0_137 (.X (dpath__PC_n_9), .A (INSTR[2]), .B (n_0_103), .S (drc_ipo_n82));
XNOR i_0_136 (.X (n_0_102), .A1 (PC[1]), .A2 (n_0_121));
MX2 i_0_135 (.X (dpath__PC_n_8), .A (INSTR[1]), .B (n_0_102), .S (drc_ipo_n82));
MX2 i_0_134 (.X (dpath__PC_n_7), .A (INSTR[0]), .B (n_0_121), .S (drc_ipo_n82));
NAND2 i_0_133 (.X (n_0_101), .A1 (INSTR[6]), .A2 (INSTR[5]));
INV4 i_0_132 (.X (n_0_100), .A (n_0_101));
NOR2 i_0_131 (.X (n_0_99), .A1 (n_0_117), .A2 (n_0_101));
    // Should become INSTR[3]
NAND2 i_0_130 (.X (n_0_98), .A1 (INSTR[3]), .A2 (n_0_100));
NOR2 i_0_129 (.X (n_0_97), .A1 (n_0_114), .A2 (drc_ipo_n79));
NOR2 i_0_128 (.X (n_0_96), .A1 (n_0_116), .A2 (n_0_115));
NAND2 i_0_127 (.X (n_0_95), .A1 (n_0_97), .A2 (drc_ipo_n84));
MX2 i_0_126 (.X (dpath_rf_n_0), .A (sgo___n_3_126), .B (\dpath_rf_rf7[3] ), .S (drc_ipo_n73));
MX2 i_0_125 (.X (dpath_rf_n_1), .A (sgo___n125), .B (\dpath_rf_rf7[2] ), .S (drc_ipo_n73));
MX2 i_0_124 (.X (dpath_rf_n_2), .A (sgo___n_2_122), .B (\dpath_rf_rf7[1] ), .S (drc_ipo_n73));
MX2 i_0_123 (.X (dpath_rf_n_3), .A (sgo___n_1_124), .B (\dpath_rf_rf7[0] ), .S (drc_ipo_n73));
NOR2 i_0_122 (.X (n_0_94), .A1 (drc_ipo_n79), .A2 (drc_ipo_n120));
NAND2 i_0_121 (.X (n_0_93), .A1 (drc_ipo_n84), .A2 (drc_ipo_n76));
MX2 i_0_120 (.X (dpath_rf_n_11), .A (sgo___n_3_126), .B (\dpath_rf_rf6[3] ), .S (drc_ipo_n109));
MX2 i_0_119 (.X (dpath_rf_n_12), .A (sgo___n125), .B (\dpath_rf_rf6[2] ), .S (drc_ipo_n109));
MX2 i_0_118 (.X (dpath_rf_n_13), .A (sgo___n_2_122), .B (\dpath_rf_rf6[1] ), .S (drc_ipo_n109));
MX2 i_0_117 (.X (dpath_rf_n_14), .A (sgo___n_1_126), .B (\dpath_rf_rf6[0] ), .S (drc_ipo_n109));
NOR2 i_0_116 (.X (n_0_92), .A1 (n_0_116), .A2 (INSTR[1]));
NOR3 i_0_115 (.X (n_0_91), .A1 (n_0_116), .A2 (n_0_114), .A3 (INSTR[1]));
NAND2 i_0_114 (.X (n_0_90), .A1 (drc_ipo_n83), .A2 (drc_ipo_n85));
MX2 i_0_113 (.X (dpath_rf_n_15), .A (drc_ipo_n114), .B (\dpath_rf_rf5[3] ), .S (drc_ipo_n80));
MX2 i_0_112 (.X (dpath_rf_n_16), .A (drc_ipo_n93), .B (drc_ipo_n98), .S (drc_ipo_n80));
MX2 i_0_111 (.X (dpath_rf_n_17), .A (sgo___n_2_122), .B (\dpath_rf_rf5[1] ), .S (drc_ipo_n80));
MX2 i_0_110 (.X (dpath_rf_n_18), .A (sgo___n_1_124), .B (drc_ipo_n97), .S (drc_ipo_n80));
NOR3 i_0_109 (.X (n_0_89), .A1 (n_0_116), .A2 (INSTR[1]), .A3 (INSTR[0]));
NAND2 i_0_108 (.X (n_0_88), .A1 (drc_ipo_n83), .A2 (drc_ipo_n86));
MX2 i_0_107 (.X (dpath_rf_n_19), .A (drc_ipo_n114), .B (drc_ipo_n96), .S (drc_ipo_n81));
MX2 i_0_106 (.X (dpath_rf_n_20), .A (drc_ipo_n93), .B (\dpath_rf_rf4[2] ), .S (drc_ipo_n81));
MX2 i_0_105 (.X (dpath_rf_n_21), .A (sgo___n_2_124), .B (\dpath_rf_rf4[1] ), .S (drc_ipo_n81));
MX2 i_0_104 (.X (dpath_rf_n_22), .A (sgo___n_1_124), .B (drc_ipo_n95), .S (drc_ipo_n81));
NOR2 i_0_103 (.X (n_0_87), .A1 (n_0_115), .A2 (INSTR[2]));
NOR4 i_0_102 (.X (n_0_86), .A1 (n_0_115), .A2 (n_0_114), .A3 (drc_ipo_n79), .A4 (INSTR[2]));
MX2 i_0_101 (.X (dpath_rf_n_23), .A (\dpath_rf_rf3[3] ), .B (sgo___n_3_126), .S (drc_ipo_n77));
MX2 i_0_100 (.X (dpath_rf_n_24), .A (\dpath_rf_rf3[2] ), .B (sgo___n127), .S (drc_ipo_n77));
MX2 i_0_99 (.X (dpath_rf_n_25), .A (\dpath_rf_rf3[1] ), .B (sgo___n_2_124), .S (drc_ipo_n77));
MX2 i_0_98 (.X (dpath_rf_n_26), .A (\dpath_rf_rf3[0] ), .B (sgo___n_1_126), .S (drc_ipo_n77));
NAND2 i_0_97 (.X (n_0_85), .A1 (drc_ipo_n76), .A2 (drc_ipo_n87));
MX2 i_0_96 (.X (dpath_rf_n_27), .A (sgo___n_3_126), .B (\dpath_rf_rf2[3] ), .S (drc_ipo_n74));
MX2 i_0_95 (.X (dpath_rf_n_28), .A (sgo___n127), .B (\dpath_rf_rf2[2] ), .S (drc_ipo_n74));
MX2 i_0_94 (.X (dpath_rf_n_29), .A (sgo___n_2_124), .B (drc_ipo_n115), .S (drc_ipo_n74));
MX2 i_0_93 (.X (dpath_rf_n_30), .A (sgo___n_1_126), .B (\dpath_rf_rf2[0] ), .S (drc_ipo_n74));
NOR2 i_0_92 (.X (n_0_84), .A1 (INSTR[2]), .A2 (INSTR[1]));
NAND2 i_0_91 (.X (n_0_83), .A1 (drc_ipo_n76), .A2 (drc_ipo_n90));
MX2 i_0_90 (.X (dpath_rf_n_31), .A (sgo___n_3_126), .B (OPORT[3]), .S (drc_ipo_n75));
MX2 i_0_89 (.X (dpath_rf_n_32), .A (sgo___n127), .B (OPORT[2]), .S (drc_ipo_n75));
MX2 i_0_88 (.X (dpath_rf_n_33), .A (sgo___n_2_124), .B (OPORT[1]), .S (drc_ipo_n75));
MX2 i_0_87 (.X (dpath_rf_n_34), .A (sgo___n_1_126), .B (OPORT[0]), .S (drc_ipo_n75));
NAND2 i_0_86 (.X (n_0_82), .A1 (n_0_120), .A2 (drc_ipo_n79));
MX2 i_0_85 (.X (n_0_81), .A (\dpath_rf_rf6[2] ), .B (\dpath_rf_rf7[2] ), .S (drc_ipo_n120));
MX2 i_0_84 (.X (n_0_80), .A (\dpath_rf_rf2[2] ), .B (\dpath_rf_rf3[2] ), .S (sgo___n122));
NAND2 i_0_83 (.X (n_0_79), .A1 (n_0_80), .A2 (drc_ipo_n87));
NAND2 i_0_82 (.X (n_0_78), .A1 (\dpath_rf_rf4[2] ), .A2 (drc_ipo_n86));
MX2 i_0_81 (.X (n_0_77), .A (OPORT[2]), .B (IPORT[2]), .S (sgo___n122));
NAND2 i_0_80 (.X (n_0_76), .A1 (n_0_77), .A2 (drc_ipo_n90));
NAND2 i_0_79 (.X (n_0_75), .A1 (drc_ipo_n98), .A2 (drc_ipo_n85));
NAND2 i_0_78 (.X (n_0_74), .A1 (n_0_79), .A2 (n_0_76));
NAND2 i_0_77 (.X (n_0_73), .A1 (n_0_78), .A2 (n_0_75));
NOR2 i_0_76 (.X (sgo__n133), .A1 (n_0_74), .A2 (n_0_73));
NAND2 i_0_75 (.X (n_0_71), .A1 (n_0_81), .A2 (drc_ipo_n84));
NAND2 i_0_74 (.X (n_0_70), .A1 (n_0_72), .A2 (n_0_71));
MX2 i_0_73 (.X (n_0_69), .A (INSTR[2]), .B (n_0_70), .S (n_0_119));
NAND2 i_0_72 (.X (n_0_68), .A1 (n_0_69), .A2 (drc_ipo_n112));
NOR2 i_0_71 (.X (n_0_67), .A1 (n_0_119), .A2 (INSTR[1]));
NAND2 i_0_70 (.X (n_0_66), .A1 (\dpath_rf_rf5[1] ), .A2 (drc_ipo_n85));
NOR2 i_0_69 (.X (n_0_65), .A1 (sgo___n122), .A2 (OPORT[1]));
NOR2 i_0_68 (.X (sgo__n131), .A1 (n_0_114), .A2 (IPORT[1]));
NOR4 i_0_67 (.X (n_0_63), .A1 (INSTR[2]), .A2 (INSTR[1]), .A3 (n_0_65), .A4 (n_0_64));
NAND2 i_0_66 (.X (n_0_62), .A1 (\dpath_rf_rf4[1] ), .A2 (drc_ipo_n86));
MX2 i_0_65 (.X (n_0_61), .A (drc_ipo_n115), .B (\dpath_rf_rf3[1] ), .S (sgo___n122));
NAND2 i_0_64 (.X (n_0_60), .A1 (n_0_61), .A2 (drc_ipo_n87));
MX2 i_0_63 (.X (n_0_59), .A (\dpath_rf_rf6[1] ), .B (\dpath_rf_rf7[1] ), .S (INSTR[0]));
NAND2 i_0_62 (.X (n_0_58), .A1 (n_0_59), .A2 (drc_ipo_n84));
NAND2 i_0_61 (.X (n_0_57), .A1 (n_0_66), .A2 (n_0_58));
NAND2 i_0_60 (.X (n_0_56), .A1 (n_0_62), .A2 (n_0_60));
NOR4 i_0_59 (.X (sgo__n_1_121), .A1 (n_0_57), .A2 (n_0_56), .A3 (INSTR[6]), .A4 (n_0_63));
NOR2 i_0_58 (.X (n_0_54), .A1 (n_0_67), .A2 (n_0_55));
NAND2 i_0_57 (.X (n_0_53), .A1 (sgo___n_2_122), .A2 (drc_ipo_n72));
MX2 i_0_56 (.X (n_0_52), .A (\dpath_rf_rf6[0] ), .B (\dpath_rf_rf7[0] ), .S (drc_ipo_n120));
NAND2 i_0_55 (.X (n_0_51), .A1 (n_0_52), .A2 (drc_ipo_n84));
NOR2 i_0_54 (.X (n_0_50), .A1 (n_0_119), .A2 (INSTR[0]));
MX2 i_0_53 (.X (n_0_49), .A (OPORT[0]), .B (IPORT[0]), .S (drc_ipo_n120));
NAND2 i_0_52 (.X (n_0_48), .A1 (n_0_49), .A2 (drc_ipo_n90));
MX2 i_0_51 (.X (n_0_47), .A (\dpath_rf_rf2[0] ), .B (\dpath_rf_rf3[0] ), .S (drc_ipo_n120));
NAND2 i_0_50 (.X (n_0_46), .A1 (n_0_47), .A2 (drc_ipo_n87));
NAND2 i_0_49 (.X (n_0_45), .A1 (n_0_48), .A2 (n_0_46));
MX2 i_0_48 (.X (n_0_44), .A (drc_ipo_n95), .B (drc_ipo_n97), .S (INSTR[0]));
NAND2 i_0_47 (.X (n_0_43), .A1 (n_0_44), .A2 (n_0_92));
NAND2 i_0_46 (.X (n_0_42), .A1 (n_0_51), .A2 (n_0_43));
NOR3 i_0_45 (.X (n_0_41), .A1 (n_0_45), .A2 (n_0_42), .A3 (INSTR[6]));
NOR2 i_0_44 (.X (n_0_40), .A1 (n_0_50), .A2 (n_0_41));
NAND2 i_0_43 (.X (n_0_39), .A1 (drc_ipo_n110), .A2 (sgo___n_1_124));
NOR2 i_0_42 (.X (n_0_38), .A1 (sgo___n_2_122), .A2 (drc_ipo_n72));
NAND2 i_0_41 (.X (n_0_37), .A1 (n_0_53), .A2 (drc_ipo_n71));
INV4 i_0_40 (.X (n_0_36), .A (n_0_37));
XNOR i_0_39 (.X (n_0_35), .A1 (sgo___n_2_122), .A2 (drc_ipo_n72));
NOR2 i_0_38 (.X (n_0_34), .A1 (slo___n191), .A2 (n_0_36));
INV4 i_0_37 (.X (n_0_33), .A (slo___n164));
NAND2 i_0_36 (.X (n_0_32), .A1 (n_0_33), .A2 (n_0_68));
NOR2 i_0_35 (.X (n_0_31), .A1 (n_0_69), .A2 (drc_ipo_n112));
NOR2 i_0_34 (.X (n_0_30), .A1 (n_0_117), .A2 (INSTR[5]));
NOR2 i_0_33 (.X (n_0_29), .A1 (n_0_118), .A2 (INSTR[3]));
NOR3 i_0_32 (.X (n_0_28), .A1 (n_0_31), .A2 (drc_ipo_n88), .A3 (drc_ipo_n89));
XNOR i_0_31 (.X (n_0_27), .A1 (drc_ipo_n112), .A2 (n_0_69));
NAND2 i_0_30 (.X (n_0_26), .A1 (n_0_32), .A2 (n_0_28));
MX2 i_0_29 (.X (n_0_25), .A (\dpath_rf_rf6[3] ), .B (\dpath_rf_rf7[3] ), .S (drc_ipo_n120));
NAND2 i_0_28 (.X (n_0_24), .A1 (n_0_25), .A2 (drc_ipo_n84));
NAND2 i_0_27 (.X (n_0_23), .A1 (\dpath_rf_rf5[3] ), .A2 (drc_ipo_n85));
MX2 i_0_26 (.X (n_0_22), .A (OPORT[3]), .B (IPORT[3]), .S (sgo___n122));
NAND2 i_0_25 (.X (n_0_21), .A1 (n_0_22), .A2 (drc_ipo_n90));
MX2 i_0_24 (.X (n_0_20), .A (\dpath_rf_rf2[3] ), .B (\dpath_rf_rf3[3] ), .S (sgo___n122));
NAND2 i_0_23 (.X (n_0_19), .A1 (n_0_20), .A2 (drc_ipo_n87));
NAND2 i_0_22 (.X (n_0_18), .A1 (drc_ipo_n96), .A2 (drc_ipo_n86));
NAND2 i_0_21 (.X (n_0_17), .A1 (n_0_21), .A2 (n_0_19));
NAND2 i_0_20 (.X (n_0_16), .A1 (n_0_23), .A2 (n_0_18));
NOR2 i_0_19 (.X (sgo__n123), .A1 (n_0_17), .A2 (n_0_16));
NAND2 i_0_18 (.X (n_0_14), .A1 (n_0_15), .A2 (n_0_24));

// Mux which drives, eventually, the accumulator
MX2 i_0_17 (.X (n_0_13), .A (INSTR[3]), .B (n_0_14), .S (n_0_119));
NOR2 i_0_16 (.X (n_0_12), .A1 (drc_ipo_n94), .A2 (drc_ipo_n88));
MX2 i_0_15 (.X (n_0_11), .A (n_0_12), .B (drc_ipo_n94), .S (n_0_13));
XOR i_0_14 (.X (n_0_10), .A1 (n_0_26), .A2 (n_0_11));
MX2 i_0_13 (.X (dpath_n_0), .A (n_0_10), .B (drc_ipo_n94), .S (drc_ipo_n78));
NOR2 i_0_12 (.X (n_0_9), .A1 (n_0_33), .A2 (drc_ipo_n89));
XNOR i_0_11 (.X (n_0_8), .A1 (n_0_27), .A2 (n_0_9));
MX2 i_0_10 (.X (n_0_7), .A (n_0_8), .B (n_0_68), .S (drc_ipo_n88));
MX2 i_0_9 (.X (dpath_n_1), .A (n_0_7), .B (drc_ipo_n112), .S (drc_ipo_n78));
NOR2 i_0_8 (.X (n_0_6), .A1 (drc_ipo_n71), .A2 (drc_ipo_n89));
XNOR i_0_7 (.X (n_0_5), .A1 (n_0_35), .A2 (n_0_6));
MX2 i_0_6 (.X (n_0_4), .A (n_0_5), .B (n_0_53), .S (drc_ipo_n88));
MX2 i_0_5 (.X (dpath_n_2), .A (n_0_4), .B (drc_ipo_n111), .S (drc_ipo_n78));
NOR2 i_0_4 (.X (n_0_3), .A1 (drc_ipo_n110), .A2 (drc_ipo_n88));
NOR2 i_0_3 (.X (n_0_2), .A1 (n_0_3), .A2 (drc_ipo_n78));
NOR2 i_0_2 (.X (n_0_1), .A1 (sgo___n_1_124), .A2 (slo___n197));
NOR2 i_0_1 (.X (n_0_0), .A1 (drc_ipo_n78), .A2 (drc_ipo_n71));
NOR2 i_0_0 (.X (dpath_n_3), .A1 (n_0_1), .A2 (n_0_0));
INV4 dpath__PC_i_3_0 (.X (dpath__PC_n_15), .A (RSTN));
DFFQ \dpath_A_reg[0]  (.Q (\dpath_A[0] ), .CLK (CLK), .D (dpath_n_3));
DFFQ \dpath_A_reg[1]  (.Q (\dpath_A[1] ), .CLK (CLK), .D (dpath_n_2));
DFFQ \dpath_A_reg[2]  (.Q (\dpath_A[2] ), .CLK (CLK), .D (dpath_n_1));
DFFQ \dpath_A_reg[3]  (.Q (\dpath_A[3] ), .CLK (CLK), .D (dpath_n_0));
DFFQ \dpath_rf_rf0_reg[0]  (.Q (drc_ipo_n102), .CLK (CLK), .D (dpath_rf_n_34));
DFFQ \dpath_rf_rf0_reg[1]  (.Q (drc_ipo_n104), .CLK (CLK), .D (dpath_rf_n_33));
DFFQ \dpath_rf_rf0_reg[2]  (.Q (drc_ipo_n106), .CLK (CLK), .D (dpath_rf_n_32));
DFFQ \dpath_rf_rf0_reg[3]  (.Q (drc_ipo_n108), .CLK (CLK), .D (dpath_rf_n_31));
DFFQ \dpath_rf_rf2_reg[0]  (.Q (\dpath_rf_rf2[0] ), .CLK (CLK), .D (dpath_rf_n_30));
DFFQ \dpath_rf_rf2_reg[1]  (.Q (\dpath_rf_rf2[1] ), .CLK (CLK), .D (dpath_rf_n_29));
DFFQ \dpath_rf_rf2_reg[2]  (.Q (\dpath_rf_rf2[2] ), .CLK (CLK), .D (dpath_rf_n_28));
DFFQ \dpath_rf_rf2_reg[3]  (.Q (\dpath_rf_rf2[3] ), .CLK (CLK), .D (dpath_rf_n_27));
DFFQ \dpath_rf_rf3_reg[0]  (.Q (\dpath_rf_rf3[0] ), .CLK (CLK), .D (dpath_rf_n_26));
DFFQ \dpath_rf_rf3_reg[1]  (.Q (\dpath_rf_rf3[1] ), .CLK (CLK), .D (dpath_rf_n_25));
DFFQ \dpath_rf_rf3_reg[2]  (.Q (\dpath_rf_rf3[2] ), .CLK (CLK), .D (dpath_rf_n_24));
DFFQ \dpath_rf_rf3_reg[3]  (.Q (\dpath_rf_rf3[3] ), .CLK (CLK), .D (dpath_rf_n_23));
DFFQ \dpath_rf_rf4_reg[0]  (.Q (\dpath_rf_rf4[0] ), .CLK (CLK), .D (dpath_rf_n_22));
DFFQ \dpath_rf_rf4_reg[1]  (.Q (\dpath_rf_rf4[1] ), .CLK (CLK), .D (dpath_rf_n_21));
DFFQ \dpath_rf_rf4_reg[2]  (.Q (\dpath_rf_rf4[2] ), .CLK (CLK), .D (dpath_rf_n_20));
DFFQ \dpath_rf_rf4_reg[3]  (.Q (\dpath_rf_rf4[3] ), .CLK (CLK), .D (dpath_rf_n_19));
DFFQ \dpath_rf_rf5_reg[0]  (.Q (\dpath_rf_rf5[0] ), .CLK (CLK), .D (dpath_rf_n_18));
DFFQ \dpath_rf_rf5_reg[1]  (.Q (\dpath_rf_rf5[1] ), .CLK (CLK), .D (dpath_rf_n_17));
DFFQ \dpath_rf_rf5_reg[2]  (.Q (\dpath_rf_rf5[2] ), .CLK (CLK), .D (dpath_rf_n_16));
DFFQ \dpath_rf_rf5_reg[3]  (.Q (\dpath_rf_rf5[3] ), .CLK (CLK), .D (dpath_rf_n_15));
DFFQ \dpath_rf_rf6_reg[0]  (.Q (\dpath_rf_rf6[0] ), .CLK (CLK), .D (dpath_rf_n_14));
DFFQ \dpath_rf_rf6_reg[1]  (.Q (\dpath_rf_rf6[1] ), .CLK (CLK), .D (dpath_rf_n_13));
DFFQ \dpath_rf_rf6_reg[2]  (.Q (\dpath_rf_rf6[2] ), .CLK (CLK), .D (dpath_rf_n_12));
DFFQ \dpath_rf_rf6_reg[3]  (.Q (\dpath_rf_rf6[3] ), .CLK (CLK), .D (dpath_rf_n_11));
DFFQ \dpath_rf_rf7_reg[0]  (.Q (\dpath_rf_rf7[0] ), .CLK (CLK), .D (dpath_rf_n_3));
DFFQ \dpath_rf_rf7_reg[1]  (.Q (\dpath_rf_rf7[1] ), .CLK (CLK), .D (dpath_rf_n_2));
DFFQ \dpath_rf_rf7_reg[2]  (.Q (\dpath_rf_rf7[2] ), .CLK (CLK), .D (dpath_rf_n_1));
DFFQ \dpath_rf_rf7_reg[3]  (.Q (\dpath_rf_rf7[3] ), .CLK (CLK), .D (dpath_rf_n_0));
DFFC \dpath__PC_PC_reg[0]  (.Q (drc_ipo_n117), .CL (dpath__PC_n_15), .CLK (CLK), .D (dpath__PC_n_7));
DFFC \dpath__PC_PC_reg[1]  (.Q (drc_ipo_n100), .CL (dpath__PC_n_15), .CLK (CLK), .D (dpath__PC_n_8));
DFFC \dpath__PC_PC_reg[2]  (.Q (slo_n214), .CL (dpath__PC_n_15), .CLK (CLK), .D (dpath__PC_n_9));
DFFC \dpath__PC_PC_reg[3]  (.Q (PC[3]), .CL (dpath__PC_n_15), .CLK (CLK), .D (dpath__PC_n_10));
DFFC \dpath__PC_PC_reg[4]  (.Q (drc_ipo_n119), .CL (dpath__PC_n_15), .CLK (CLK), .D (dpath__PC_n_11));
DFFC \dpath__PC_PC_reg[5]  (.Q (PC[5]), .CL (dpath__PC_n_15), .CLK (CLK), .D (dpath__PC_n_12));
DFFC \dpath__PC_PC_reg[6]  (.Q (PC[6]), .CL (dpath__PC_n_15), .CLK (CLK), .D (dpath__PC_n_13));
BUF4 drc_ipo_c77 (.X (drc_ipo_n87), .A (slo___n232));
BUF4 drc_ipo_c86 (.X (drc_ipo_n96), .A (\dpath_rf_rf4[3] ));
BUF4 drc_ipo_c84 (.X (drc_ipo_n94), .A (\dpath_A[3] ));
BUF4 drc_ipo_c80 (.X (drc_ipo_n90), .A (n_0_84));
BUF4 drc_ipo_c85 (.X (drc_ipo_n95), .A (\dpath_rf_rf4[0] ));
BUF4 drc_ipo_c81 (.X (drc_ipo_n91), .A (\dpath_A[0] ));
BUF4 drc_ipo_c78 (.X (drc_ipo_n88), .A (slo___n224));
BUF4 drc_ipo_c88 (.X (drc_ipo_n98), .A (\dpath_rf_rf5[2] ));
BUF4 drc_ipo_c83 (.X (drc_ipo_n93), .A (\dpath_A[2] ));
BUF4 drc_ipo_c90 (.X (OPORT[0]), .A (drc_ipo_n102));
BUF4 drc_ipo_c89 (.X (PC[1]), .A (drc_ipo_n100));
BUF4 drc_ipo_c87 (.X (drc_ipo_n97), .A (\dpath_rf_rf5[0] ));
BUF4 drc_ipo_c82 (.X (drc_ipo_n92), .A (\dpath_A[1] ));
BUF4 drc_ipo_c76 (.X (drc_ipo_n86), .A (n_0_89));
BUF4 drc_ipo_c75 (.X (drc_ipo_n85), .A (n_0_91));
BUF4 drc_ipo_c79 (.X (drc_ipo_n89), .A (n_0_29));
BUF4 drc_ipo_c74 (.X (drc_ipo_n84), .A (n_0_96));
BUF4 drc_ipo_c73 (.X (drc_ipo_n83), .A (n_0_99));
BUF4 drc_ipo_c72 (.X (drc_ipo_n82), .A (n_0_113));
BUF4 drc_ipo_c71 (.X (drc_ipo_n81), .A (n_0_88));
BUF4 drc_ipo_c70 (.X (drc_ipo_n80), .A (n_0_90));
BUF4 drc_ipo_c69 (.X (drc_ipo_n79), .A (n_0_98));
BUF4 drc_ipo_c68 (.X (drc_ipo_n78), .A (n_0_82));
BUF4 drc_ipo_c67 (.X (drc_ipo_n77), .A (n_0_86));
BUF4 drc_ipo_c66 (.X (drc_ipo_n76), .A (slo___n150));
BUF4 drc_ipo_c65 (.X (drc_ipo_n75), .A (n_0_83));
BUF4 drc_ipo_c64 (.X (drc_ipo_n74), .A (n_0_85));
BUF4 drc_ipo_c63 (.X (drc_ipo_n73), .A (n_0_95));
BUF4 drc_ipo_c62 (.X (drc_ipo_n72), .A (n_0_54));
BUF4 drc_ipo_c61 (.X (drc_ipo_n71), .A (n_0_39));
BUF4 drc_ipo_c91 (.X (OPORT[1]), .A (drc_ipo_n104));
BUF4 drc_ipo_c92 (.X (OPORT[2]), .A (drc_ipo_n106));
BUF4 drc_ipo_c93 (.X (OPORT[3]), .A (drc_ipo_n108));
BUF4 drc_ipo_c94 (.X (drc_ipo_n109), .A (n_0_93));
BUF4 drc_ipo_c95 (.X (drc_ipo_n110), .A (n_0_40));
BUF4 drc_ipo_c96 (.X (drc_ipo_n111), .A (drc_ipo_n92));
BUF4 drc_ipo_c97 (.X (drc_ipo_n112), .A (drc_ipo_n93));
BUF4 drc_ipo_c98 (.X (drc_ipo_n113), .A (drc_ipo_n91));
BUF4 drc_ipo_c99 (.X (drc_ipo_n114), .A (drc_ipo_n94));
BUF4 drc_ipo_c100 (.X (drc_ipo_n115), .A (\dpath_rf_rf2[1] ));
BUF4 drc_ipo_c101 (.X (PC[0]), .A (drc_ipo_n117));
BUF4 drc_ipo_c102 (.X (PC[4]), .A (drc_ipo_n119));
BUF4 drc_ipo_c103 (.X (drc_ipo_n120), .A (INSTR[0]));
INV4 sgo___L1_c104 (.X (sgo___n121), .A (drc_ipo_n120));
INV4 sgo___L2_c105 (.X (sgo___n122), .A (sgo___n121));
BUF4 sgo__c106 (.X (n_0_15), .A (sgo__n123));
INV4 sgo___L1_c107 (.X (sgo___n124), .A (drc_ipo_n112));
INV4 sgo___L2_c108 (.X (sgo___n125), .A (sgo___n124));
INV4 sgo___L3_c109 (.X (sgo___n126), .A (sgo___n125));
INV4 sgo___L4_c110 (.X (sgo___n127), .A (sgo___n126));
INV1 sgo___L1_c_3_104 (.X (sgo___n_3_121), .A (n_0_111));
INV4 sgo___L2_c_3_105 (.X (sgo___n_3_122), .A (sgo___n_3_121));
INV4 sgo___L1_c_3_108 (.X (sgo___n_3_125), .A (drc_ipo_n114));
INV4 sgo___L2_c_3_109 (.X (sgo___n_3_126), .A (sgo___n_3_125));
INV4 sgo___L1_c_2_104 (.X (sgo___n_2_121), .A (drc_ipo_n111));
INV4 sgo___L2_c_2_105 (.X (sgo___n_2_122), .A (sgo___n_2_121));
INV4 sgo___L3_c_2_106 (.X (sgo___n_2_123), .A (sgo___n_2_122));
INV4 sgo___L4_c_2_107 (.X (sgo___n_2_124), .A (sgo___n_2_123));
BUF4 sgo__c_1_104 (.X (n_0_55), .A (sgo__n_1_121));
INV4 sgo___L1_c_1_106 (.X (sgo___n_1_123), .A (drc_ipo_n113));
INV4 sgo___L2_c_1_107 (.X (sgo___n_1_124), .A (sgo___n_1_123));
INV4 sgo___L3_c_1_108 (.X (sgo___n_1_125), .A (sgo___n_1_124));
INV4 sgo___L4_c_1_109 (.X (sgo___n_1_126), .A (sgo___n_1_125));
BUF4 sgo__c114 (.X (n_0_64), .A (sgo__n131));
BUF4 sgo__c116 (.X (n_0_72), .A (sgo__n133));
INV1 slo___L1_c118 (.X (slo___n135), .A (n_0_104));
INV4 slo___L2_c119 (.X (slo___n136), .A (slo___n135));
INV1 slo___L1_c124 (.X (slo___n141), .A (n_0_106));
INV4 slo___L2_c125 (.X (slo___n142), .A (slo___n141));
INV4 slo___L1_c132 (.X (slo___n149), .A (n_0_94));
INV1 slo___L2_c133 (.X (slo___n150), .A (slo___n149));
INV4 slo___L1_c146 (.X (slo___n163), .A (n_0_34));
INV4 slo___L2_c147 (.X (slo___n164), .A (slo___n163));
INV1 slo___L1_c173 (.X (slo___n190), .A (n_0_38));
INV4 slo___L2_c174 (.X (slo___n191), .A (slo___n190));
INV1 slo___L1_c179 (.X (slo___n196), .A (n_0_2));
INV4 slo___L2_c180 (.X (slo___n197), .A (slo___n196));
INV1 slo___L1_c187 (.X (slo___n204), .A (slo_n214));
INV4 slo___L2_c188 (.X (PC[2]), .A (slo___n204));
INV4 slo___L1_c193 (.X (slo___n215), .A (n_0_107));
INV4 slo___L2_c194 (.X (slo___n216), .A (slo___n215));
INV1 slo___L1_c201 (.X (slo___n223), .A (n_0_30));
INV4 slo___L2_c202 (.X (slo___n224), .A (slo___n223));
INV1 slo___L1_c209 (.X (slo___n231), .A (n_0_87));
INV4 slo___L2_c210 (.X (slo___n232), .A (slo___n231));

endmodule //core


